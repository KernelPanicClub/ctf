BZh91AY&SY�o �߀Py����߰?���Py����@�i�& i��dhш�F� �@sbh0�2d��`�i���!�H�"�FFLM�~��� ���SA�	���dɓ#	�i�F& �"BhF��L�Sh�( Ѡ2=&j$��AED+��% f��楤���/�ga�D�,Ж���6�V+Z����~�S��,Sj���e�w���B�ޥ,�>橳��n#��6�ls�I�v�Mpkw �Ca�IzFc|k���,Y���!"�ʓI �ąo��u��iP-6G;݄дxK�D920eא1M_��g�\�$�:��l.N�W��e�l�����7�V�]ַ��[�E},jE�2��nn	�[{��WW8+k�T��������7���m��Sp��~"$��?%l�YȘ!�DP�cK�v��m[ť�0����B����$[H1�֏�2����j��xyG��x�z��|\�a���ք�'�	��K� Uc�v����WL�����:�4�e����5l�G������lc��6"���΄kk�4)�)|�9��g�A?06��9�����IB��CN�J�h2���2:�ZA0t�J�9d�g&H�"rSD����V��'�&�h	�����뜂�D�iz�1A�9�鈛2S��vi�Z;J.�X��C
�J�����w�_ >f��i膔��dP����L{�� 6�b�!���4;��Y�C0|�����IXQw���4lY0G��w�r7���(�]���� �a0ța��SC����d��,)B�x���6�$-{$� �+��)4u�%!���t���܃���/��e(����y*�,�:�:̈���߸�bI���\R�cK��?Ñ�3�ζ���
�k&6)?<�:�f>���o�u������Nb�!C+m�-�F�,�Á�^b&,��C5�;	�����
����ijX��r ��J�R1	�A����|'{b����e��Qt�	."	�
����)���x`